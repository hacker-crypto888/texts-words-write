b0VIM 7.4      ���]|  $  root                                    kmaster                                 ~root/upload_web_app/src/index.js                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            utf-8U3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      s            U   t         h   �         ~   1     	   J   �     
   \   �        �   U        �   �        J   ^        N   �        P   �        �   F        \   �        n   ,        a   �        ]   �        V   X           �        @   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ad  .        s   �  �  �  �  X  0  �  �  �  [     �  �    X  $     �  �  n  H    �  �  �  Z  -  �
  �
  �
  z
  V
  *
  �	  �	  z	  P	  9	  '	  	  �  �  �  �  �  �  y  d  S  9  )      �  �  �  �  �  �  f  P  6      �  �  �  �  �  v  b  H  *      �  �  �  �  �  �  h  R  K  G  /  �  �  v  4    �  �  �  �  �  �  s  e  O  B  :  6  5    �  �  �  �  �  �  �  j  N                                                    if(document.getElementById('myAudioFiles').hasChildNodes) {     event.preventDefault();   disableButton = (event) => {      }     this.btn.removeAttribute("disabled");     event.preventDefault();   handleWordInput = (event) => {   }     event.preventDefault();   handleSubmit = (event) => {    }     });         null       wordinputError:         null,       audioplayerToggle:     this.setState({   fieldOnblur = () => {    }     dataOutput.appendChild(someData);     someData.id = 'some-data';     const someData = document.createElement('a');     const dataOutput = document.getElementById("outputJsonFile");     const allAudioElements = document.getElementsByTagName('audio');      this.btn.setAttribute('disabled','disabled');      document.getElementById('loadingAudioFiles').hidden = true;   componentDidMount() {   }     };       firstAudio:null       myAudioItems:null,       someData:null,       dataOutput:null,       dataLists:null,       allAudioElements:null,       idx:null,       element:null,       myarray:null,       indexes:[],       previewAudioFiles:null,       audioElements:null,       preview:null,       previewMyItems:null,       myAudioNode:null,       itemsImportMode:null,       wordInputField:null,       myAudioFiles:null,       myBlub:null,       myBlob:null,       sourceFile:null,       theFirstChild:null,       sourceTag:null,       audioFilePreview:null,       myAudio:null,       audioId:null,       mp3WordList:null,       audioplayerToggle:"",       user: '',       emailError:'',       nameError:'',       email: '',       name: '',       wordinputError: '',       items: [],       controls:true,       mountElements:[],       variableErrors:'',       targetValue: '',       checkTarget:'',       wordtest:'',       checkInput:'',       inputValue:'',     this.state = {     super(props);   constructor(props) { class BasicForm extends React.Component { document.head.appendChild(s);  s.onload = function(e){ /* now that its loaded, do something */ };  s.src = "https://cdnjs.cloudflare.com/ajax/libs/jquery/3.4.1/jquery.min.js"; const s = document.createElement("script"); const mammoth = require("mammoth"); //const textract = require('textract'); //const officeParser = require('officeparser'); //const dxe = require('docx-extractor'); //const anyFileParser = require('anyfileparser'); //const docxParser = require('docx-parser'); //  generateHtml = office2html.generateHtml; //const office2html = require('office2html'), //const docxParser = require('docx-parser'); //const WordExtractor = require("word-extractor"); //const converter = require('office-converter')(); //const unoconv = require('unoconv'); //const getDocumentProperties = require('office-document-properties'); //const word2html = require('word2html'); //const docx = require('./docx') //const pdf = require('pdf-parse'); //const PdfReader = require("pdfreader").PdfReader; //const pdfText = require('pdf-text'); //pdfjsLib.workerSrc = pdfjsWorkerBlobURL; //const pdfjsWorkerBlobURL = URL.createObjectURL(pdfjsWorkerBlob); //const pdfjsWorkerBlob = new Blob([pdfjsWorker]); //const PDFExtract = require('pdf.js-extract').PDFExtract; //const pdfjsWorker = require('pdfjs-dist/build/pdf.worker.min'); const fs = require('fs'); const path = require('path'); pdfjsLib.GlobalWorkerOptions.workerSrc = '//mozilla.github.io/pdf.js/build/pdf.worker.js'; const pdfjsLib = require('pdfjs-dist'); import DatePicker from 'react-date-picker'; import axios from 'axios'; import './index.css'; import ReactDOM from 'react-dom';  import React, {setState} from 'react';  ad  �  �     @   �  �  �  �  }  h  !     �  �  i  W  $      �  �  �  �  �  �  �  t  �  �  �  �    �  �  �  E  "    �
  �
  �
  -
  $
  �	  �	  �	  �	  �	  �	  1	  
	  �  �  �  y  x    �  a  7  6  4  &          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ReactDOM.render(<BasicForm />, document.getElementById('root'));  }   }     );       </form>            <div id={`download_zone`}></div>          <div id={`download_all_items`}></div>          <a id={`download_items`} ref={a => {this.a = a}} onClick={this.downloadItems} download={`items.json`} href={``} ></a>         <input type={`submit`} value={`Submit entered text`} className={`btn btn-success btn-block`} />            </button>           Add a new text         <button onClick={this.addNewText} className={`btn btn-success btn-block`}>           </label>           {this.state.textareaIsEmpty}           <br /><textarea onChange={this.handleTextChange} placeholder="Enter a text" value={this.state.value} />             Your Text:         <label id={`labelText`}>          <pre id={`display`}></pre>         <div id={`outputpdf`}></div>                  <iframe id={`processor`} src={`http://hubgit.github.com/2011/11/pdftotext/`}></iframe>         <iframe id={`input`} type={`application/pdf`} />         <p id={`result3`}></p>         <p id={`result2`}></p>         <p id={`result1`}></p>         <div id={`preview`}></div>   	<div id={`dropzone`} multiple onDragEnter={this.onDragEnter} onDrop={this.onDrop} onDragOver={this.onDragOver}></div>          </div>           <label for="subscribeNews">I have no database.json</label>           <input type="checkbox" id={`noDatabaseFile`} value={this.state.noDatabaseFile} onChange={this.checkBox} />         <div>         </div>           <label for="playAllTheWords">Play all the words</label>           <input type="checkbox" id="playAllTheWords" value={this.state.preloadOrAutoplay} onChange={this.checkBox} name="playAllTheWords"/>         <div>       <form enctype={`multipart/form-data`} onSubmit={this.handleSubmittedText}>     return (       }       }, true);         //};           }             break;               //console.log(event.data.cleanup());               //}               //   return this.toLowerCase().replace(/[^a-zA-Z0-9]+/g, "-").split('-');               //String.prototype.cleanup = function() {               console.log(event.data);                outputpdf.textContent = event.data.replace(/\s+/g, " ");             default:             // anything else = the processor has returned the text of the PDF                    break;                xhr.send(); ad  �  !        �  �  _  X  9  �  �  �  �  i  9    �  p  2  !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           };                 //console.log(JSON.stringify(this.response));                 //console.log(processor.contentWindow.postMessage(this.response, "*"));                 processor.contentWindow.postMessage(this.response, "*");               xhr.onload = (event) => {               xhr.responseType = "arraybuffer";               xhr.open('GET', input.getAttribute("src"), true);                const xhr = new XMLHttpRequest;             case "ready":             // "ready" = the processor is ready, so fetch the PDF file           switch (event.data){                  if (event.source !== processor.contentWindow) return;         //window.onload = (event) => {       window.addEventListener("message", function(event){ ad  .  �     V   U  0    �  �  �  �  �  �  �  e  ^  �  |  `  N  B  *      �  �  �  M  C  ;  5  4  �  �  �  �  �  G    �
  �
  �
  �
  ~
  <
  5
  1
  
  �  �  p  U  F  <     �  �  �  p  j  f  L  !  �  �  �  �  �  �  �  s  _  R  7  /  �  �    y  @    �  �    {  n  L    �  �  �  l  T  (  '  �  �  �  N  �  �  �  �                           };               //console.log(JSON.stringify(this.response));               //console.log(processor.contentWindow.postMessage(this.response, "*"));               processor.contentWindow.postMessage(this.response, "*");             xhr.onload = (event) => {             xhr.responseType = "arraybuffer";             xhr.open('GET', input.getAttribute("src"), true);              const xhr = new XMLHttpRequest;           case "ready":           // "ready" = the processor is ready,      const outputpdf = document.getElementById("outputpdf");       const processor = document.getElementById("processor");       const input = document.getElementById('input');     if (processor && input.src) {   render() {   }     console.log(event.currentTarget.value);      console.log(this.state.value);      console.log(importedTexts.dataset.textValue);      console.log(document.getElementById('wordinput').value);     importedTexts.dataset.textValue += this.state.value;     }       importedTexts.dataset.textValue = "";     if(importedTexts.dataset.textValue ===(null||undefined||false)) {     const importedTexts = document.getElementById('preview');     });         event.target.value       value:     this.setState({   addNewText = (event) => {   }      }       myElements[0].play();     if (myElements && myElements.length) {      const myElements = document.getElementsByTagName('audio');     //const allAudioElements = this.state;   autoplay = (event) => {   }     }       document.getElementById('noDatabaseFile').removeAttribute('checked');        } else {       //this.handleText();       document.getElementById('dropzone').hidden = true;       console.log("alert");       });           true         jsonSecondConfirm:       this.setState({       document.getElementById('noDatabaseFile').checked = true;     if (/*this.state.value.replace(/[!?:;.,]+/g, "").replace(/(\r\n|\n|\r)/gm,"") !== "" &&*/ document.getElementById('noDatabaseFile').checked === false && document.getElementById('preview').innerHTML === "" && window.confirm("You dropped no file. Ok to continue and generate a new database or Cancel and upload a file.")) {   alertNoDatabaseFile = (event) => {   }     }        //document.getElementById('noDatabaseFile').checked = true;       document.getElementById('dropzone').hidden = true;       });           true          jsonSecondConfirm:        this.setState({     } else if (document.getElementById('noDatabaseFile').checked) {       document.getElementById('dropzone').hidden = false;       });           false         jsonSecondConfirm:        this.setState({     if (!document.getElementById('noDatabaseFile').checked && this.state.jsonSecondConfirm === true) {      }       }         }           droppedFiles.removeChild(droppedFiles.firstChild);           while (droppedFiles.hasChildNodes()) {         const droppedFiles = document.getElementById('preview');         });             []           myItems:         this.setState({         });             false           databaseIsLoaded:         this.setState({       if (this.state.databaseIsLoaded === true && window.confirm("the database is to be removed. To remove the database anyway, press ok. Press cancel to keep your database loaded in the dropzone.")) {              console.log("checkbox");     if (document.getElementById('noDatabaseFile').checked) {      }       }         }           el.currentTime = 0;           el.pause();         el.onended = (event) => {       for (let el of audioTagName) {     if (!document.getElementById('playAllTheWords').checked && audioTagName && audioTagName.length && Object.keys(audioTagName)[0].onended !== (null||undefined||false)) { ad     z     U   �  �  N  *    �  �  �  }  H  3  �  �  �  �  �  �  �  �  �  �  p  8        �  �  �  l  f  I  H  �  �  �    \  �
  �
  �
  8
  
  �	  �	  m	  &	  �  �  �  s  ?    �  �  �  1  �  �  �  <  �  �  �  �  v    �  �  �  R  �  �  q  p  �  �        �  �  �  �  z  y                              ////const mylist = ['a', 'b', 'a', 'c', 'a', 'd'];               //const indexes = [];             }               };                 }                    //myAudioItems.insertBefore(event.currentTarget, myAudioItems.children[indexAudioElement]);                   myAudioItems.childNodes[indexAudioElement].play();                   //event.currentTarget.remove();                   const indexAudioElement = Array.prototype.indexOf.call(myAudioItems.children, event.currentTarget) + 1;                    //const firstAudio = allAudioElements[0];                   const myAudioItems = document.getElementById('myAudioFiles');                   //const allAudioElements = document.getElementsByTagName('audio');                   //allAudioElements[0].play();                   //allAudioElements[0].remove();                    //oItems.firstChild.play();                   //myAudioItems.appendChild(firstAudio);                   //const myAudioItems = document.getElementById('myAudioFiles');                          //allAudioElements[0].remove();                      //const firstAudio = allAudioElements[0];                   //const allAudioElements = document.getElementsByTagName('audio');                 if (allAudioElements && allAudioElements.length && allAudioElements.length >= 2) {                 //if (allAudioElements[1]) {                 //allAudioElements[0].remove();                  //console.log(event.currentTarget);                 const allAudioElements = document.getElementsByTagName('audio');               audioFilePreview.onended = (event) => {             if (document.getElementById('playAllTheWords').checked) {             }               event.currentTarget.currentTime = 0;             audioFilePreview.onpause = (event) => {             audioFilePreview.controls=true;             audioFilePreview.id=item.word;             audioFilePreview.key=item.id;             audioFilePreview.className=item.word;             const audioFilePreview = document.createElement('audio');              //const myAudioFiles = document.getElementById('myAudioFiles');             //console.log(item);           items.forEach(function(item, index, object) {           const items = myBlub.items;           const myBlub = JSON.parse(document.getElementById('items_by_date').dataset.databaseJson);           document.getElementById('loadingAudioFiles').hidden = false;          if(document.getElementById('items_by_date') && document.getElementById('items_by_date').dataset.databaseJson) {       .then(function(mp3WordList){       })         return response.json();       .then(function(response){     fetch("https://raw.githubusercontent.com/nathanielove/English-words-pronunciation-mp3-audio-download/master/ultimate.json")      const myAudioFiles = [];     }       myNode.removeChild(myNode.firstChild);     while(myNode.firstChild) {     const myNode = document.getElementById('myAudioFiles');   displayAudio = event => {   };     });       this.validateName();     this.setState({ name: event.target.value }, () => {   handleNameChange = event => {   }     });         ''        controls:      this.setState({   disableFormButton = () => {   }     }       });           targetValue === '' ? 'play a word' : null         checkTarget:           inputValue === '' ? 'enter a word' : null,         checkInput:           inputValue === targetValue ? this.removeAudioPlayer() : null,               wordtest:       this.setState({       //console.log({inputValue});       //console.log({targetValue});       this.btn.setAttribute("disabled", "disabled");       const { inputValue } = this.state;       const targetValue = document.getElementById('wordinput').dataset.targetValue; ad     �     h   �  �  e  A    �  �  �  �  �  �  �  X    �  �  �  6  �  �  h  !  �  �  �  b        �
  �
  ~
  n
  ^
  Q
  	
  
  �	  �	  �	  f	  4	  (	  	  	  �  �  �  �  h  A  -    �  �  �  y  U  A  +  �  �  �  �  b  1  +      �  �  �  �  �  �  �  �  w  v  u     �  �  �  �  /    �  �  �  [  -  �  �  �  j  R  ;  :  (  '  �  �  �                     Start a new game                <button id={`loadItemsForNewGame`} onClick={this.displayAudio}>             </div>               </button>                click me              <button ref={btn => { this.btn = btn; }} onClick={this.disableButton} >              />                                onChange={e => this.setState({ inputValue: e.target.value }) }                onFocus={this.handleWordInput}                onClick={this.handleWordInput}                //onMouseOver={this.displayAudio}                value={this.state.inputValue}                placeholder='Enter word'                id={`wordinput`}                className={`form-control ${this.state.wordinputError ? 'is-invalid' : ''}`}              <input              <label htmlFor={`wordinput`}></label>              </div>                <span className="sr-only">Loading...</span>              <div className="spinner-border" id={`loadingAudioFiles`} role="status">              <div className={`form-group`}>        <form onSubmit={this.handleSubmit}>     return(        render() {       }     });         ''       inputValue:     this.setState({     }       mountElements.removeAttribute('controls');       mountElements.currentTime = 0;       mountElements.pause();     if (mountElements !== undefined) {     });         mountElements === undefined ? "Please choose and listen to a word first" : null       variableErrors:     this.setState({     //console.log({mountElements});     const mountElements = document.getElementById(targetValue);     //console.log({targetValue});     });         `Values: \n ${inputValue} / ${targetValue} ok`          wordtest:     this.setState({     const { inputValue } = this.state;     const targetValue = document.getElementById('wordinput').dataset.targetValue;   removeAudioPlayer = (props) => {   }      //display AUDIO FILES THAT ARE IN AN ARRAY ONE BY ONE          })         });           previewMyAudioFiles.appendChild(item);          myAudioFiles.forEach(function(item, index, object) {         const previewMyAudioFiles = document.getElementById('myAudioFiles');         }           });              document.getElementById('loadingAudioFiles').hidden = true;                          });               }                                  myAudioFiles.push(audioFilePreview);                 //myAudioFiles.appendChild(audioFilePreview);                 })                    audioFilePreview.insertBefore(sourceFile, theFirstChild);                   sourceFile.type = 'audio/mpeg';                    sourceFile.className = item.word;                    //console.log(mp3link);                   sourceFile.src = mp3link;                    const sourceFile = document.createElement('source');                   const theFirstChild = audioFilePreview.firstChild;                 mp3[1].forEach(function(mp3link, indexmp3link, objectmp3link) {               if(mp3[0] === item.word && mp3[1].length){             [...Object.entries(mp3WordList)].forEach(function(mp3, indexmp3, objectmp3) {             //console.log(item.word);             };               wordInputField.dataset.targetValue = audioFilePreview.id;               const wordInputField = document.getElementById('wordinput');             audioFilePreview.onplay = (event) => {                                              //console.log(indexes);               //}               //  idx = mylist.indexOf(element, idx + 1);               //  indexes.push(idx);               //while (idx != -1) {               //const idx = mylist.indexOf(element);               //const element = event.currentTarget;               //const mylist = allAudioElements; ad  Q   ]     ~   �  �  �  �  z  K    �  �  �  ;      �  �  �  {  V  A    �  �  �  �  �  �  �  �  �  `  I  8  %    �  �  �  �  �  �  �  |  g  T  =  *    �
  �
  �
  �
  �
  �
  
  k
  Q
  6
   
  
  �	  �	  �	  �	  �	  �	  x	  h	  T	  @	  +	  	  		  �  �  �  �  �  �  �  �  c  K  4      �  �  �  �  �  x  ^  C  .        �  �  �  |  C    �  �  F    �  �  r  L  H  /    �  �  �  z  8    �  �  �  �  �  ]  \                                                                                   if(document.getElementById("download_items").dataset.databaseJson.length) {    handleSubmittedDate = (event) => {   }     }       myInputNode.removeChild(myInputNode.firstChild);     while(myInputNode.firstChild) {     const myInputNode = document.getElementById('inputJsonFile');     //}     //  myNode.removeChild(myNode.firstChild);     //while(myNode.firstChild) {     //const myNode = document.getElementById('outputJsonFile');     this.setState({ date });   onChange = (date) => {   }     dataOutput.appendChild(someData);     someData.id = 'some-data';     const someData = document.createElement('a');     const dataOutput = document.getElementById("outputJsonFile");     document.getElementById('dropzoneSortByDate').hidden = true;     document.getElementById('submit-date-btn').hidden = true;     document.getElementById('labelJsonInPublicDir').hidden = true;     document.getElementById('jsonInPublicDir').hidden = true;     document.getElementById('labelDropMyJson').hidden = true;     document.getElementById('dropMyJson').hidden = true;     document.getElementById('dropzoneSortByDate').hidden = false;     this.setState({date});     const date = new Date();   componentDidMount() {   }     }       dataOutput:null       someData:null,       myDatabaseJson:null,       myPreviewNode:null,       myOutputNode:null,       myInputNode:null,       myNode:null,       downloadLink:null,       downloadAll:null,       jsonString:null,       saveFile:null,       importMode:null,           noFileType:null,       myItems:null,           databaseIsLoaded:null,       myBlub:null,       myBlob:null,       thirdres:null,       response:null,       fd:null,       k:null,       j:null,       i:null,       dt:null,       reader:null,       fileName:null,       preview:null,       myImage:null,       img:null,       file:null,        files:null,       outputLink:null,       outputJson:null,       addLink:'',       content:"",       mydatepicker:null,       listContents:null,       jsonContent:"",       allItemsByDate:null,       myItemsByDate:null,       myItems:null,       jsonString:null,       myNewBlob:null,       element:null,       res:null,       mynewDb:null,       downloadLink:null,       daysDate:new Date(),       today:null,       myBlub:null,       myDatabase:null,       myBlob:null,       response:null,       valueArray:null,       url:null,       text:null,       shortArray:'',       json:null,       data:null,       database:[],       selectedDate:'',       date: '',     this.state = {     super(props)   constructor(props) { class FillInTheDateForm extends React.Component {  }   }     );           </form>            </div>             </div>               </div>                 <FillInTheDateForm />               <div id={`myFillInTheDateForm`}>               </div>                 <RegistrationForm />               <div>             <div className="card card-body">            <div className="collapse" id="mysettings">            </p>              </button>               {`\u2699`} Settings              <button class="btn btn-primary" type="button" data-toggle="collapse" data-target="#mysettings" aria-expanded="false" aria-controls="collapseExample">            <p>             <div id={`myAudioFiles`}></div>            <div>{this.state.variableErrors}</div>            <div>{this.state.checkTarget}</div>            <div>{this.state.checkInput}</div>            <div>{this.state.wordtest}</div>               <br />              </button> ad     O     J   �  �  �  z  �  �  �  �  h  9    	  �  �  �  �  �  p  E  �  �  �  �  �  _  ^      �  �  �  Y  3  �
  
  �	  �	  S	  	  	  �  [  /    �  �  �  ,      �  �  �  z  7    �  �  �  d  �  �    �  r  0  �  A     �  �  �  �  O  N                         //const myOutputNode = document.getElementById('outputJsonFile');         //INITIALIZE DOWNLOAD LINKS AREA//       } else {          outputJson.appendChild(outputLink);         //COLUMNS: WORD, ID, ARRAY OF DATES (PROGRAM JAVASCRIPT)         outputLink.dataset.databaseJson = JSON.stringify({"items": myItemsByDate}); //LINES: UNKNOWN         //WHERE THE DATABASES (IN CONSTANTS) ARE LOADED / ASSIGNED: LOOK FOR ITS LINES AND COLUMNS IN THE CODE ABOVE IT (USING THE PROPS)         //////////////------------------------------------------/         //EVENT LISTENERS CAN ONLY BE WORKED OUT IF THE JSON IS CORRECTLY WORKED OUT AS WELL         //////////////------------------------------------------/         //BOOTSTRAP\\\\\\ CAN ONLY BE POSSIBLE IF ALL THE INFO FROM FETCH (FROM THE DROPPED FILES) AND THE BLOBS (DATABASES THAT ARE MADE WITH THE FORMDATA) IS COMPLETE         //////////////------------------------------------------/         //DATA INPUT(FOR THE AUDIO DISPLAYER)/OUTPUT(FOR THE FORM FIELDS) TO DISPLAY AUDIO IS A DATASET         //////////////------------------------------------------/         //2)DATASET          //STORE IN: 1) JSON         //////////////------------------------------------------/         //FILE TYPES (FETCH)          //ARRAYS / OBJECTS FIELDS (EX: NAME, WORD, ID, DATE, TITLE         //ARRAY TYPES / OBJECTS TYPES         //DATASET TYPES         //BLOB TYPE         //////////////------------------------------------------/          //DATASET TYPE: JSON         //alert('Your JSON file with items sorted by date is ready. save it under public/ directory of your app, reload page and start playing!');         outputJson.hidden = false;          outputLink.hidden = false;         outputLink.id = 'items_by_date';         outputLink.download = 'items.json';         outputLink.innerHTML = "download JSON file (date of data entry: "+selectedDate+ ")";         //\\THE DATASET WAS ASSIGNED TO ITS HTML ELEMENT ELSEWHERE IN THE CODE          //DATE OF EACH WORD (SEVERAL DATES FOR SEVERAL DAYS OF OCCURRENCE)         //IT WAS NOT PRECISED WHETHER DATA CAME FROM A FILE WITH SOME TYPE OR JUST THE TEXT TYPED IN THE TEXT AREA         //COLUMNS: WORD, ID, DATES OF CONSULTATION         //ORIGIN: DATASET          outputLink.href = URL.createObjectURL(new Blob([JSON.stringify({"items": [...myItemsByDate]},null,2)], {type: 'application/json'})); //OBJECT TYPE: ARRAY         //BLOB TYPE: JSON, \\\\\\NO MORE NEEDED (THE APP CAN DIRECTLY LOAD THE WORDS THAT WERE DROPPED IN THE DROPZONE//////         //console.log(myItemsByDate);         const outputLink = document.createElement('a');         }           document.getElementById("items_by_date").remove();         if(document.getElementById("items_by_date")) {                  const outputJson = document.getElementById("outputJsonFile");          //CREATES OUTPUT JSON FILE DOWNLOAD LINK           }           myInputNode.removeChild(myInputNode.firstChild);         while(myInputNode.firstChild) {         const myInputNode = document.getElementById('inputJsonFile');         //INITIALIZE DOWNLOAD LINKS AREA//       if ([...myItemsByDate].length){        //  //FROM THERE, THE ARRAY "MY ITEMS BY DATE" IS USED TO OUTPUT THE DOWNLOAD LINk            });         }                      myItemsByDate.push(item);          if(item.dates.includes(selectedDate)){       myItems.items.forEach(function(item, index, object) {       console.log(myItems);        const myItemsByDate = [];       //console.log(myItems);       const selectedDate = (this.state.date.getMonth()+1)+'/'+this.state.date.getDate()+'/'+this.state.date.getFullYear();         //MY DATE PICKER                  const myItems = JSON.parse(document.getElementById("download_items").dataset.databaseJson); ad     �     \   �  �  �  D    �  �  �  �  g  1  �  �  �  b  ?      �  �  �  �  �  �  �  v    �  �  �  9  	    �
  u
  t
  (
  �	  �	  S	  	  �  �  �  �  �  �  �  P  (  �  ~     �  b  U  N  �  �  �  }  a  >    �  �  �  �  M  @    �  �  �  �  �  �  �  �  y  f  V  E  �  �  �  l  8    �  �  �     I must advance the colours of my love Perforce, against all cheques, rebukes and manners, In such a righteous fashion as I do, Good Mistress Page, for that I love your daughter than I can: you may ask your father; here he comes. his dole! They can tell you how things go better motions: if it be my luck, so; if not, happy man be with you. Your father and my uncle hath made       value: '',/*`Truly, for mine own part, I would little or nothing       email: '',       name: '',     this.state = {     super(props);   constructor(props) { class RegistrationForm extends React.Component {  }   }       );       </form>       <div id={`outputJsonFile`}></div>       <div id={`inputJsonFile`}></div>       </div>         <input type="submit" id="submit-date-btn" value="Submit selected date" className='btn btn-success btn-block' />         <div>       </div>         />           value={this.state.date}           onMouseOver={this.itemsByDateLoadForm}           onChange={this.onChange}           id="myDatePicker"         <DatePicker       <div>       <div id={`previewSortByDate`}></div>       <div id={`dropzoneSortByDate`} multiple onDragEnter={this.onDragEnter} onDrop={this.onDrop} onDragOver={this.onDragOver}></div>              </div>         <label id={`labelDropMyJson`} for={`dropMyJson`}> Rather load my own database.json file</label>         <input type={`radio`} id={`dropMyJson`} value={`drop`} name={`importMode`} />         <label id={`labelJsonInPublicDir`} for={`jsonInPublicDir`}>Sort items by date</label>         <input type={`radio`} id={`jsonInPublicDir`} value={`load`} name={`importMode`} />       <div id={`setImportMode`} onChange={event => this.setImportMode(event)}>       <label>Load words by date</label>       <form onSubmit={this.handleSubmittedDate}>     return (       render() {       }     }                //document.getElementById('dropzoneSortByDate').removeAttribute('hidden');       document.getElementById('submit-date-btn').removeAttribute('hidden');       document.getElementById('labelJsonInPublicDir').removeAttribute('hidden');       document.getElementById('jsonInPublicDir').checked = true;       document.getElementById('dropzoneSortByDate').hidden = true;       document.getElementById('jsonInPublicDir').removeAttribute('hidden');        document.getElementById('labelDropMyJson').removeAttribute('hidden');       document.getElementById('dropMyJson').removeAttribute('hidden');        //console.log(event.target.clientHeight);       event.target.removeEventListener('mouseover', this.itemsByDateLoadForm);        }         document.getElementById("items_by_date").remove();       if(document.getElementById("items_by_date")) {     if (document.getElementById('items_by_date') && document.getElementById('items_by_date').dataset.databaseJson) {     //alert('test');   itemsByDateLoadForm = (event) => {   }      }                //=====/=/=/=/=/=/=/=/=/=/=/=/=/         //=====/=/=/=/=/=/=/=/=/=/=/=/=/       }         outputJson.hidden = false;         outputLink.hidden = false;         outputJson.appendChild(outputLink);         outputLink.id = 'noitem';         outputLink.textContent = 'no item corresponds to your request.';         const outputLink = document.createElement('p');         const someData = document.createElement('a');         const outputJson = document.getElementById("outputJsonFile");         //OUTPUTS TEXT FOR NO VALID ITEM          }           myInputNode.removeChild(myInputNode.firstChild);         while(myInputNode.firstChild) {         const myInputNode = document.getElementById('inputJsonFile');         //}         //  myOutputNode.removeChild(myOutputNode.firstChild);         //while(myOutputNode.firstChild) { ad     K     �   �  �    P  +  �  �  �  �  T    �  �  �  S         �  �  �  �  �  �  y  i  Z  I  ;  -    �  �  �  �  �  �  u  `  Q  B  2     
  �
  �
  �
  �
  �
  u
  _
  S
  E
  /
   
  
  �	  �	  �	  �	  �	  �	  �	  i	  N	  /	  	  �  �  �  �  t  V  <  %    �  �  �  �  �  c  Q  5      �  �  �  �  �  d  K  4      �  �  �  �  l  V  B  ,    �  �  �  �  �  �  m  O  8  $    �  �  �  �  �  �  q  Z  C  &  	  �  �  �  �  �  �  �  w  _  K  J                       pdfUtil:null,       arrayBuffer:null,       reader:null,       xhr:null,       loadFile:null,       absPath:null,       path:null,       fs:null,       messages:null,       html:null,       thisIsMyWordList:null,       thisIsMyTextList:null,       allMyTexts:null,       allMyWords:null,       myTextId:null,       myTextList:null,       myResult:null,       c:null,       allMyTexts:null,       result:null,       myBiggestWordList:null,       mySuperWordList:null,       newText:null,       myWordInfo:null,       allWordsFromTexts:null,       myTextContent:null,       output:null,       finalArray:null,       myTextInfo:null,       importedTexts:null,       newTexts: null,       myDivForNewData:null,       mySuperList:null,       indataset:null,       newText:null,       jsonParse:null,       msTime:Date.now(),       allTheImportedTexts:null,       contentOfThisText:null,       infoAboutThisText:null,       allTheImportedTexts:null,       daysDate:null,       indexAudioElement:null,       firstAudio:null,       audioTagName:null,       preloadOrAutoplay:null,       someData:null,       dataOutput:null,       indexCurrentAudio:null,       allElementsButOne:null,       myElements:null,       aNewHtmlElement:null,       aNewElement:null,       myItemsFromText:null,       items:null,       myDatabaseForUpload:null,       itemsWereDropped:null,       textareaIsEmpty:null,       textAtFileCreation:null,       databaseJson:null,       downloadLink:null,       downloadAll:null,       allMyItems:null,       wordsFromText:null,       wordsFromDatabase:null,       compilationOfWordsFromDatabase:null,       previewMyDatabase:null,       compilationOfWordsFromText:null,       mapJson:null,       droppedFiles:null,       databaseIsLoaded:false,       jsonSecondConfirm:false,       daysDate:new Date(),       noDatabaseFile:false,       fileName:null,       noFileType:null,       myImage:null,       myBlob:null,       myBlub:null,       img:null,       preview:null,       file:null,       dt:null,       emailError: '',       a:null,       x:[],       wordIdItems:[],       wordIdKVPairs:new Set(),       testdatabase:[],       newItem:null,       jsonItemsMap:new Map(),       wordsIdMap:new Map(),       arrays:[],       duplicate:null,       items:null,       map:null,       n: null,       m: null,       loadedText:[],       datesFromDatabase:[],       wordList:[],       downloadArray:[],       concatArray:null,       nameError: '',       bigDatabase:[],       itemlist:"",       databaseLength:null,       l:null,       k:null,       concat:[],       word:{},       today:'',       j:null,       database:[],       textError:'',       blobData:[],       date:new Date(),       itemList:[],       importText:'',       text:'',       i:null, my two mistresses: what a beast am I to slack it!`,*/ I must of another errand to Sir John Falstaff from as my word; but speciously for Master Fenton. Well, three; for so I have promised, and I'll be as good Fenton had her; I will do what I can for them all Master Slender had her; or, in sooth, I would Master would my master had Mistress Anne; or I would fire and water for such a kind heart. But yet I A kind heart he hath: a woman would run through Her father will be angry. Till then farewell, sir: she must needs go in; And as I find her, so am I affected. My daughter will I question how she loves you, I will not be your friend nor enemy: Come, trouble not yourself. Good Master Fenton, And not retire: let me have your good will. ad  0   D     �   �  �  �  �  �  �  r  b  N  >  .      �  �  �  �  �  �  ~  k  [  G  6  #       �  �  �  �  �  w  a  H  2  +  $  #  �  �  �  �  �  �  O  +  �  �  ]  >    �
  �
  W
  >
  #
  
  �	  �	  �	  �	  �	  �	  �	  �	  �	  |	  D	  )	  !	  	  	  �  �  �  �  �  �  ~  ]  I  8  �  �  �  �  �  �  �  �  4  ,  (    �  �  �  l  `  \  C    �  �  �  �  �  �  �  �  O    �  �  �  I      �  �  4  ,  +    �  e  D  C                                                  const daysDate = new Date();     //YOU IMPORT THE TEXT YOU ENTERED INTO THE VARIABLE WORDLIST     //if (/*this.state.value.replace(/[!?:;.,]+/g, "").replace(/(\r\n|\n|\r)/gm,"") === ""*/) {     //ALERT BOXES (TEXT IN TEXTAREA)      //}     //if (document.getElementById('noDatabaseFile').checked === true && this.state.myItems === ([]||undefined)) {     console.log(importedTexts.dataset.textValue);     //importedTexts.dataset.textValue += this.state.value;     //}     //  importedTexts.dataset.textValue = "";     //if (importedTexts.dataset.textValue === undefined) {     const importedTexts = document.getElementById('preview');     //}     //  this.state.value = document.getElementById('preview').dataset.textValue;     //if (this.state.value === (null||undefined)) {     //YOU HAVE NO DATABASE.JSON AND YOU HAVE NO ITEMS     //const wordList = [];   handleText = (event) => {    }            //const importText = importedTexts.dataset.splitContent;     const importedTexts = document.getElementById('preview');   splitContent = () => {   }     //  });     //    this.setState({ database });     //    const database = res.data.items.map(obj => obj);     //  .then(res => {     //axios.get(`./database.json`)   importAllWords = (event) => {   }     });         email.length > 3 ? null : 'Email must be longer than 3 characters'        emailError:     this.setState({     const { email } = this.state;   validateEmail = () => {    }     });         name.length > 3 ? null : 'Name must be longer than 3 characters'       nameError:     this.setState({     const { name } = this.state;   validateName = () => {    };     });       this.validateEmail();     this.setState({ email: event.target.value }, () => {   handleEmailChange = event => {    };     });       this.validateName();     this.setState({ name: event.target.value }, () => {   handleNameChange = event => {    }         //allTheImportedTexts = {};     const allMyTexts = [];      const thisIsMyTextList = [];     const thisIsMyWordList = [];     const allMyWords = [];     const wordList = [];     importedTexts.dataset.textValue = '';     const importedTexts = document.getElementById('preview');     //const allTheImportedTexts = document.getElementById('preview').dataset.textImport;     dataOutput.appendChild(someData);     someData.id = 'some-data';     const someData = document.createElement('a');     const dataOutput = document.getElementById("outputJsonFile");     document.getElementById('noDatabaseFile').addEventListener('checked', this.checkBox);     this.a.removeAttribute("href");     window.addEventListener('drop',this.windowdrop);     window.addEventListener('dragover',this.windowdragover);   componentDidMount() {    }      this.handleSubmittedText = this.handleSubmittedText.bind(this);      };              pdfAsArray:null       pdfAsDataUri:null,       rawLength:null,       raw:null,       base64:null,       base64Index:null,       BASE64_MARKER:null,       returnedBase64:null,       returnedBlob:null,       img:null,       binary:null,       base64:null,       text:null,       display:null,       arr:null,       length:null,       bloburl:null,       blob:null,       m:null,       dataurl:null,       outputpdf:null,       processor:null,       input:null,       options:null,       pdfExtract:null,       arr:null,       enc:null,       bufView:null,       buf:null,       pdffile3:null,       pdffile2:null,       pdffile1:null,       rows:null,       pdfBuffer:null,       myFile:null,       pdf_path:null, ad  
   F     J   �  �  �  �  �  y    �  �  B    �  h  a  D  $    �  U  '  �
  �
  �
  c
  1
  �	  �	  �	  �	  [	  -	  ,	  �  �  �  �  �  X  8  �  |  b  X  C    �  �  }  `  =    [  �  (  '  &  %  $  #  �  �  �  �    �  V    �  �  �  �  �  R  F  E                //}         //  importedTexts.dataset.words = [];         //if (importedTexts.dataset.words === (undefined||null)) {          }           mytext.pop();           //console.log(mytext);           //console.log(importedTexts.dataset.splitContent); //String in Array           importedTexts.dataset.splitContent = mytext[6][1]; //importedTexts.dataset.splitContent IS A STRING THAT CONTAINS THE TEXTUAL CONTENT OF THE FILE           //console.log(mytext[6][1]);         if (mytext && mytext.length === 7){ //mytext IS AN OBJECT THAT CONTAINS INFO ABOUT THE TEXT OF THE FILE         //json word by word          //}         //  importedTexts.dataset.words = [];          //if(importedTexts.dataset.words === (undefined||null)) {              const myTextId = Math.random().toString(16).substring(7); //myTextIf IS A STRING THAT WAS GENERATED RANDOMLY BY THE PROGRAM AS A TEXT ID TO RECOGNIZE WHICH WORD BELONGS TO WHICH TEXT AND CONVERSELY       allMyTexts.forEach(function(mytext) { //mytext IS A JSON ARRAY THAT CONTAINS INFO ABOUT A TEXT       const allMyTexts = JSON.parse(importedTexts.dataset.texts); //allMyTexts is a JSON ARRAY THAT CONTAINS ALL THE TEXTS HAVING BEEN INSERTED, DROPPED OR ADDED TO BE HANDLED BY THE PROGRAM       const thisIsMyTextList = [];       const thisIsMyWordList = [];       const myTextList = [];     if(importedTexts.dataset.texts && JSON.parse(importedTexts.dataset.texts).length) {     //TO HAVE DROPPED FILES     //const wordList = [];     //////////////////////////////////////////////////     // - export JSON     // -      //- import PDF, DOC,      ///////////////////////////////////////////////////     //else if you imported JSON and texts OR if you imported texts and did not import JSON(add JSON import at the end of else loop)     //if you only imported JSON     ///////////////////////////////////////////////////     //const databaseJson = [];     //const importText = '';     //console.log(allTheImportedTexts);          //console.log(this.state.allTheImportedTexts);      //const allTheImportedTexts = this.state;     //indataset.push(Object.entries(newText).map(([k,v]) => [k,v]));     //const indataset = Object.entries(allTheImportedTexts).map(([k,v]) => [k,v]);      //}     //  //importedTexts.dataset.texts.push(newText);     //  console.log(importedTexts.dataset.texts);     //if(importedTexts.dataset.texts && importedTexts.dataset.texts.length) {     }       //console.log(JSON.parse(importedTexts.dataset.texts));       //console.log(importedTexts.dataset.texts);       //importedTexts.dataset.textValue = "";       importedTexts.dataset.texts = [JSON.stringify(myTextInfo.map(Object.entries))];       //importedTexts.dataset.texts = [JSON.stringify(myTextInfo.map(Object.entries))];       //console.log(myTextInfo);       myTextInfo.push(newText);       const myTextInfo = [];            } else if (importedTexts.dataset.texts === (null||undefined) && importedTexts.dataset.textValue !== "") {       //console.log(JSON.parse(importedTexts.dataset.texts));       //importedTexts.dataset.textValue = "";       importedTexts.dataset.texts=JSON.stringify([...JSON.parse(importedTexts.dataset.texts), myTextInfo.map(Object.entries)[0]]);       myTextInfo.push(newText);       const myTextInfo = [];     if (importedTexts.dataset.texts && importedTexts.dataset.texts.length && importedTexts.dataset.textValue !== "") {     //TO HAVE IMPORTED TEXTS     const mySuperList = this.state;     const newText = {"lastModified": this.state.msTime, "lastModifiedDate":this.state.today, "name": "", "webkitRelativePath": "", "size": "", "type": "", "mycontent":importedTexts.dataset.textValue};      const msTime = Date.now();     const today = (daysDate.getMonth()+1)+'/'+daysDate.getDate()+'/'+daysDate.getFullYear(); ad  9   �     N   �  �  I  j  6  �  �  �  c  +  �  �  "     �  �  �  �     �
  �
  U
  ,
  	
  �	  �	  v	  ;	  :	  �  �  �    B  �  �  %  $  �  �  �  �  �  �  �  �  [  G  !    �  �  �       �  �  �  �  �  v  N  3    �  �  �  n  Q  E  +    �  �  �  �  �  �  �                                                              //  if (b.word === "") { return; }        //  console.log(b.lastModified);       //  console.log(b);       });         console.log(a);         console.log(b);         myResult.push(a);         });           a[data[0]]=data[1]         b.forEach(function(data){         const a = {};          //console.log()       result.forEach(function(b) { //result is a JSON OBJECT THAT CONTAINS WORD AND INFO       console.log(result);       const myResult = [];       //console.log(myBiggestWordList);       //});       //        //  myBiggestWordList.push(a);       //  });       //    a[data[0]]=data[1]       //  output.forEach(function(data){       //  const a = {};        //const mySuperWordList = JSON.parse(importedTexts.dataset.wordList).forEach(function(output) {       //const wordList = this.state;       //const result = [];        const result = JSON.parse(importedTexts.dataset.wordList);       const output = [];       //const myBiggestWordList = [];       //Text import       console.log(JSON.parse(importedTexts.dataset.wordList));       });          }           });                             }             //  console.log(JSON.parse(importedTexts.dataset.wordList));                importedTexts.dataset.wordList = [JSON.stringify(myWordInfo.map(Object.entries))];             } else if (myWordInfo !== (null||undefined) && importedTexts.dataset.wordList === (null||undefined)) {               //console.log(JSON.parse(importedTexts.dataset.wordList));               //console.log(importedTexts.dataset.wordList);               //console.log(JSON.parse(importedTexts.dataset.wordList));                importedTexts.dataset.wordList = JSON.stringify([...JSON.parse(importedTexts.dataset.wordList), myWordInfo.map(Object.entries)[0]]); //importedTexts.dataset.wordList IS A JSON STRING THAT CONTAINS THE WORD LIST OF THE FORM THAT WAS JUST SUBMITTED             if (myWordInfo !== (null||undefined) && importedTexts.dataset.wordList !== (null||undefined)) {              //console.log(importedTexts.dataset.wordList);             //console.log(myWordInfo);             myWordInfo.push(output);             const myWordInfo = []; //myWordInfo IS AN ARRAY OF OBJECTS             //console.log(output);             output['myTextId']=myTextId;             output["word"]=word; // output is AN OBJECT THAT CONTAINS THE PRINCIPAL INFO ABOUT THE WORD AND ITS TEXT             });               output[data[0]]=data[1]             mytext.forEach(function(data){ //mytext IS A JSON ARRAY THAT CONTAINS ALL THE INFORMATION ABOUT THE TEXT THAT WAS DROPPED OR CREATED             const output = {};               if (word === "") { return; }              //console.log(mytext);              //console.log(word);            importedTexts.dataset.words.split(',').forEach(function(word) { //importedTexts.dataset.words IS AN ARRAY OF STRINGS THAT ARE THE WORDS OF THE TEXT THAT HAS BEEN SPLITTED INTO STRINGS OF WORDS            //console.log(importedTexts.dataset.mywords.type);           //console.log(importedTexts.dataset.mywords);           //importedTexts.dataset.mywords = importedTexts.dataset.words.split(',');           });             //console.log(importedTexts.dataset.words);             //importedTexts.dataset.words.push(element);             return (element !== (null||undefined));           importedTexts.dataset.words = x(importedTexts.dataset.splitContent.split(/[\s.?:;!,]+/)).map(function(y){ return y.replace(/[\W_]+/g," ") }).map(function(x){ return x.toLowerCase() }).filter(function( element ) {         if(importedTexts.dataset.splitContent !== (null||undefined)) {         const x = (list) => list.filter((v,i) => list.indexOf(v) === i);         //const wordList = this.state; ad     U     P   B  !  �  �  �  c  7    �  �  �  �  �  x  I  +    �  �  _  5    �  �  �  �  v  l  M  &    �
  �
  p
  '
  &
  �	  �	  �	  r	  /	  �  �  c  <    �  �  �  �  q    �  �  �  �  �  t  '  �  �  �  �  �  �  O  D  �  �  �  5  
  �  �  U      �  �  U           //const myTest = this[b.word].texts.some(v => v === myTextInfo.map(Object.entries)[0]);           //}          //for (var i=0; i<this[b.word].texts.length ; i++) {         //}         //  this[b.word].texts.push(myTextInfo.map(Object.entries)[0]);         //if(!this[b.word].texts.includes(myTextInfo.map(Object.entries)[0])) {         //console.log(myTextInfo.map(Object.entries)[0]);         //console.log(this[b.word].texts);         //console.log(this[b.word].texts);         //this[b.word].texts = JSON.stringify([...JSON.parse(this[b.word].texts), myTextInfo.map(Object.entries)[0]]);          //} else if(this[a.word].texts && this[a.word].length > 0){         //  this[a.word].texts = [JSON.stringify(myTextInfo.map(Object.entries))];         //         //if(this[a.word].texts && this[a.word].length === 0) {         //}             //}           //importedTexts.dataset.result = [Object.entries(this[b.word])];           //  importedTexts.dataset.result = [];           //} else if (importedTexts.dataset.result === (null||undefined)) {             //importedTexts.dataset.result = [...importedTexts.dataset.result, this[b.word]];           //if (importedTexts.dataset.result !== (null||undefined) && importedTexts.dataset.result && importedTexts.dataset.result.length && importedTexts.dataset.result.length > 0) {              //--------------------------------------------------------       //console.log(JSON.parse(importedTexts.dataset.addedTexts));       //importedTexts.dataset.bigTextList = JSON.stringify(myTextList.map(Object.entries));       }, Object.create(null));         }           thisIsMyTextList.push(this[f.myTextId]);            this[f.myTextId] = JSON.stringify(myTextList.map(Object.entries));         if (!this[f.myTextId]) {       myTextList.forEach(function(f) {       //importedTexts.dataset.addedTexts = JSON.stringify(myTextList.map(Object.entries));       //--------------------------------------------------------       //importedTexts.dataset.bigWordList = '';       //console.log(JSON.parse(importedTexts.dataset.addedWords));       //importedTexts.dataset.bigWordList = JSON.stringify(output.map(Object.entries));       }, Object.create(null));         }           thisIsMyWordList.push(this[f.myTextId]);            this[f.myTextId] = JSON.stringify(output.map(Object.entries));         if (!this[f.myTextId]) {       output.forEach(function(f) {       //importedTexts.dataset.addedWords = JSON.stringify(output.map(Object.entries));       console.log(output);       //const myTextList = this.state;       }, Object.create(null));         }           myTextList.push(myTextInfo);                  if (myTest === false) {         console.log(myTextList.length);         console.log(myTest);         console.log(myTextInfo.myTextId);         console.log(myTextList.myTextId);         const myTest = myTextList.some(v => v.myTextId === myTextInfo.myTextId);         //myTextInfo["myTextId"] = f.myTextId;         //delete myTextInfo[f.myTextId];         delete myTextInfo["word"];         const myTextInfo = f;         this[f.word].textsId.push(f.myTextId);         const myTextId = this.state;         //textId         }           output.push(this[f.word]);            this[f.word] = { "word": f.word, "textsId": [] };         if (!this[f.word]) {         importedTexts.dataset.wordInfo = f;         //const myTextList = this.state;       myResult.forEach(function(f) {       console.log(myResult); //OBJECT CONTAINS LIST OF WORDS AND THEIR INFO       //  myTextInfo.push(newText);       //  const myTextInfo = [];       //  const newText = {"lastModified": b.lastModified, "lastModifiedDate": b.lastModifiedDate, "name": b.name, "webkitRelativePath": b.webkitRelativePath, "size":b.size, "type":b.type}; ad     [     �   �  �  �  �  s  e  d        �  �  �  �  �  �  [  Z  S  4    �  �  �  �  �  u    �  �  �  �  �  |  t  s  Z  7  �  �  �  �  �  �  �  R  -  &  �
  �
  �
  �
  �
  �
  ^
  Y
  X
  S
  R
  /
  .
  -
  
  �	  �	  b	  Z	  4	  	  	  �  �  �  �  �  V  L  F  B  A  "      �  �  D    �  �  �  �  �  �  �  q  U  Q  P  3    �  �  �  �  �  �  �  y  _  C  (  "          �  �  �  �  �  u  S  1    �  �  �  ~  ]  Q     �  �  �  �  �  [  Z                                       if (file.name.slice(-4) === ".ods") {            }             this.sendDocxFile(file);           if (file.name.slice(-5) === ".docx") {            }             this.sendTextFile(file);           if (file.name.slice(-4) === ".txt") {            }             this.sendFile(file);           if (file.name === "database.json") {            const file = files[i];       for (let i=0; i<files.length; i++) {       //===JSON UPLOAD===//       this.dropbox(files);       console.log(files[0].name);       console.log(files[0].type);       const files = dt.files;     if(dt.files.length) {  		const dt = event.dataTransfer; 		event.preventDefault(); 		event.stopPropagation();   onDrop = (event) => {     }     } 			event.preventDefault(); 			event.stopPropagation();     if(dt.files.length) { 		const dt = event.dataTransfer;   onDragOver = (event) => {    }     } 			event.preventDefault(); 			event.stopPropagation();     if(dt.files.length) { 		const dt = event.dataTransfer;   onDragEnter = (event) => {    }     event.preventDefault();   windowdragover = (event) => {    }     event.preventDefault();   windowdrop = (event) => {    }      document.getElementById('download_items').href = url;     const url = window.URL.createObjectURL(blobData);     const blobData = new Blob([JSON.stringify({"items": this.state.wordIdItems},null,2)], {type: 'application/json'});     console.log(this.state.wordIdItems);   downloadItems = (event) => {   }     this.setState({date});   handleDateChange = date => {    }     }       });           "The text input field is empty. You cannot proceed."         textareaIsEmpty:       this.setState({     } else {       this.handleText();     if(this.state.value !== null) {      }       this.a.textContent = "";       this.a.removeAttribute('href');       }         document.getElementById('databaseAfterNewText').remove();       if(document.getElementById('databaseAfterNewText')) {     if(this.state.textAtFileCreation !== null) {     event.preventDefault();     handleSubmittedText = event => {    }            //console.log(importedTexts.dataset.result.length);     //console.log(importedTexts.dataset.result);                //button to add several texts       //remove duplicate array: no duplicate text                //console.log(this[a.word]);         //importedTexts.dataset.result.push(this[a.word]);                //importedTexts.dataset.result.push(this[a.word]);      //}     //const today = (daysDate.getMonth()+1)+'/'+daysDate.getDate()+'/'+daysDate.getFullYear();     //const daysDate = new Date();     //UPDATES DAY'S DATE      });         this.state.value       textAtFileCreation:     this.setState({      //this.a.setAttribute("href","items.json");       //ACTIVATION OF ONE DOWNLOAD LINK     //if(document.getElementById('noDatabaseFile').checked && this.state.value !== "") {     //YOU HAVE NO DATABASE.JSON AND YOU ENTERED A TEXT       }       this.alertNoDatabaseFile();     if (document.getElementById('noDatabaseFile').checked === false) {     result.length = 0;     const result = this.state;     };        //importedTexts.dataset.result = JSON.stringify(result);       //console.log(result);         //}, Object.create(null));         //}          //console.log(this[b.word].texts);                     //this[b.word].texts.push(myTextInfo.map(Object.entries)[0]);          //});           //}            //  return;           //if(text === myTextInfo.map(Object.entries)[0]) {         //{         //console.log(myTest); ad     �     \   �  �  �  {  n  b  Z  :  4  0    �  �  �  �  o  f  D  $  �  �  �  �  �  \  �  �  3  )           �
  �
  �
  T
  P
  O
  6
  
  �	  �	  �	  �	  �	  j	  =	  	  �  �  �  �  }  K  )    �  �  �  h  �  �  K  3      �  �  �  �  �  �  s  J  !    �  �  a  
  �  �  �  �  �  8  	  �  �  �  �  �                  console.log(newText);         const newText = {"lastModified": file.lastModified, "lastModifiedDate":file.lastModifiedDate, "name": file.name, "webkitRelativePath": file.webkitRelativePath, "size": file.size, "type": file.type, "mycontent":resultObject.value};         const importedTexts = document.getElementById('preview');         //console.log(resultObject.value)         result2.innerHTML = resultObject.value       mammoth.extractRawText({arrayBuffer: arrayBuffer}).then(function (resultObject) {        console.timeEnd();       })         console.log(resultObject.value)         result1.innerHTML = resultObject.value       mammoth.convertToHtml({arrayBuffer: arrayBuffer}).then(function (resultObject) {       const result3 = document.getElementById('result3');       const result2 = document.getElementById('result2');       const result1 = document.getElementById('result1');       // debugger       const arrayBuffer = reader.result;     reader.onloadend = function(event) {     const reader = new FileReader();     console.time();   sendDocxFile = (file) => {   }     console.log(this.state.myBlob);       })         });             true           databaseIsLoaded:         this.setState({         document.getElementById('noDatabaseFile').removeAttribute('checked');         document.getElementById('preview').appendChild(myDatabaseForUpload);         myDatabaseForUpload.dataset.databaseJson = JSON.stringify({"items":[...Object.entries(myItems).map(([k, v]) => [k,v])]});         myDatabaseForUpload.href = "";         myDatabaseForUpload.id = "items_by_date";                  const myDatabaseForUpload = document.createElement('a');         console.log(myItems);         this.setState({myItems});         const myItems = thirdres.map(obj => obj);       .then(thirdres => {       })         return myBlob;         console.log(file.name);         console.log(myBlob); //database.json         const myBlob = [...Object.values(myBlub.items)];         console.log(myBlub); //database.json       .then(function(myBlub) {       })         return response.json();       .then(function(response) {     fetch(URL.createObjectURL(file))     fd.append('myFile', file);     const fd = new FormData();   sendFile = (file) => {    }         //array of arrays containing columns: text imported, file type, file name, text content,         //text FILE         //this.handleText();             //this.handleText(value);                           })         }           importedTexts.dataset.texts = [JSON.stringify(myTextInfo.map(Object.entries))];         } else if (importedTexts.dataset.texts === (null||undefined)) {           importedTexts.dataset.texts=JSON.stringify([...JSON.parse(importedTexts.dataset.texts), myTextInfo.map(Object.entries)[0]]);         if (importedTexts.dataset.texts !== (null||undefined)) {         myTextInfo.push(newText);         const myTextInfo = [];         console.log(newText);         const newText = {"lastModified": file.lastModified, "lastModifiedDate":file.lastModifiedDate, "name": file.name, "webkitRelativePath": file.webkitRelativePath, "size": file.size, "type": file.type, "mycontent":valueText};         const importedTexts = document.getElementById('preview');         console.log(valueText);       .then(function(valueText) {       })         return response.text();       .then(function(response) {     fetch(URL.createObjectURL(file))     fd.append('myFile', file);     const fd = new FormData();   sendTextFile = (file) => {   }     }       //===END JSON UPLOAD===//       }           }                          this.sendPdfFile(file);           if (file.name.slice(-4) === ".pdf") {            }             this.sendOdsFile(file); ad     �     n   �  �  ~  �  �  U  K  B  ;          �  �  �  �  v  :  �  �  �  �  �  c  8      �  �  �  �  h  @  8  7    �
  �
  �
  �
  �
  R
  
  �	  �	  �	  �	  U	  	  �  �  �  c  I  #  �  �  �  �  �  �  S  +  !    �  �  �  �  }  L  *  �  �  �  �  }  7  
  �  �  �  k  I  *      �  �  �  b  X  W  Q  1    �  �  �  �  �  �  �  �  A  $  #  �  �            //  console.log(pdf);       //pdfjsLib.getDocument(arr).then(function(pdf) {        //buf.onload = () => {       //console.log(JSON.stringify(btoa(buf.split('base64,')[1])));       //console.log(JSON.stringify(btoa(atob(buf.split('base64,')[1]))));          //console.log(atob(base64));     //console.log(base64);     //const base64 = this.state;     reader.readAsDataURL(file);     }        //}       //  //input.addEventListener('load', () => URL.revokeObjectURL(URL.createObjectURL(file)), {once: true});       //  //URL.createObjectURL(file);        }         input.src = url;       } else {         input.srcObject = url;       if ('srcObject' in input) {       log('Fetching with ajax...');       log('Blob URL is: ' + url);       log('Inserting an img...');       log('Created a png blob of size: ' + blob.size);       const url = URL.createObjectURL(blob);       const blob = new Blob([pdfAsArray], {type: 'application/pdf'});       //console.log(pdfAsDataUri.isArray());       //console.log(pdfAsArray.isArray());        //}       //  return String.fromCharCode.apply(null, new Uint8Array(buffer));       //function ab2str(buffer) {       //const binary = fixBinary(atob(base64));        const pdfAsArray = convertDataURIToBinary(pdfAsDataUri);               //console.log(pdfAsDataUri);       }         return array;         console.log(array);         }           array[i] = raw.charCodeAt(i);         for(var i = 0; i < rawLength; i++) {                          console.log(array);         //const array = new ArrayBuffer(rawLength);         const array = new Uint8Array(new ArrayBuffer(rawLength));         const rawLength = raw.length;         console.log(raw);         const raw = window.atob(base64);         console.log(base64);         const base64 = dataURI.substring(base64Index);         console.log(base64Index);         const base64Index = dataURI.indexOf(BASE64_MARKER) + BASE64_MARKER.length;       function convertDataURIToBinary(dataURI) {              const BASE64_MARKER = ';base64,';       console.log(pdfAsDataUri[0].type);       const pdfAsDataUri = reader.result;       //const base64 = JSON.stringify(reader.result.split('base64,')[1]);       //const base64 = JSON.stringify(ab2str(reader.result));               //const buf = new Uint8Array(reader.result);       //console.log(reader.result);     reader.onloadend = (file) => {     const reader = new FileReader();      }         display.innerHTML += "\n" + text;     function log(text) {     display.innerHTML = (display.innerHTML || '');     const display = document.getElementById('display');     //}     //  return buf;     //  }     //    arr[i] = bin.charCodeAt(i);     //  for (var i = 0; i < length; i++) {     //  const arr = new Uint8Array(buf);     //  const buf = new ArrayBuffer(length);     //  const length = bin.length;     //function fixBinary (bin) {      const outputpdf = document.getElementById("outputpdf");     const processor = document.getElementById("processor");     const input = document.getElementById('input');   sendPdfFile = (file) => { //https://github.com/brianc/node-pdf-text   }    sendOdsFile = (file) => {    }      reader.readAsArrayBuffer(file);     };       })         }           importedTexts.dataset.texts = [JSON.stringify(myTextInfo.map(Object.entries))];         } else if (importedTexts.dataset.texts === (null||undefined)) {           importedTexts.dataset.texts=JSON.stringify([...JSON.parse(importedTexts.dataset.texts), myTextInfo.map(Object.entries)[0]]);         if (importedTexts.dataset.texts !== (null||undefined)) {         myTextInfo.push(newText);         const myTextInfo = []; ad     �     a   �  �  �  �  v  Z  !  �  �  �  �  �  �  x  .    �  �  �  ~  v  u  S  ,    �  �  �  c  b  &  �  �  �  �  e  ,  	  �
  �
  f
  
  �	  �	  o	  S	  ;	  	  �  �  �  �  �  �  <    �  �  ~  r  h  B  A    �  �  �  �  s  J    �  �    J  -    �  �  �  �  H    �  �  y  L    �  �  �  �  x  a  D    �  �                      //    .sort((y1, y2) => parseFloat(y1) - parseFloat(y2)) // sort float positions     //  Object.keys(rows) // => array of y-positions (type: float)     //function printRows() {     //const rows = {};     //});       //});         //if (item.text) console.log(item.text);         //else if (!item) callback();         //if (err) callback(err);       //new PdfReader().parseBuffer(pdfBuffer, function(err, item) {       // pdfBuffer contains the file content     //fs.readFile(pdfBuffer.name, (err, pdfBuffer) => {     //pdfBuffer.readAsArrayBuffer(file);     //const pdfBuffer = URL.createObjectURL(file);      //const result3 = document.getElementById('result3');     //const result2 = document.getElementById('result2');     //const result1 = document.getElementById('result1');     //const reader = new FileReader();     //});     //    console.log(item.text);     //  if(item && item.text)     //, function(err, item){     //console.log(pdffile3.readAsText(file).result);     //const pdffile3 = new FileReader();     //console.log(pdffile2.readAsArrayBuffer(file).result);     //const pdffile2 = new FileReader();     //console.log(pdffile1.readAsBinaryString(file).result);     //const pdffile1 = new FileReader();     //console.log(file);     //new PdfReader().parseFileItems(     //const reader = new FileReader();     //URL.createObjectURL      //reader.readAsBinaryString(file);     //reader.readAsArrayBuffer(file);      //reader.readAsArrayBuffer(file);     //});       //});       //  console.log(chunks.join(' '));        //pdfText(reader.result, function(err, chunks) {       // blob sous la forme d'un tableau typé       // reader.result contient le contenu du       //console.log(enc.readAsBinaryString(new Blob([new Uint8Array(buf)])));        //}       //    });       //        });       //            console.log(pages);       //            return pages.join("\r\n");       //        })).then(function(pages) {       //            });       //                });       //                    }).join(' ');       //                        return item.str;       //                    return textContent.items.map(function(item) {       //                return page.getTextContent().then(function(textContent) {       //            return pdf.getPage(pageNumber + 1).then(function(page) {       //        return Promise.all(pages.map(function(pageNumber) {       //        }       //            pages.push(i);       //        for (var i = 0; i < pdf.numPages; i++) {       //        var pages = [];       //    return PDFJS.getDocument(buf).then(function(pdf) {        //    pdfjsLib.cMapPacked = true;       //    pdfjsLib.cMapUrl = 'js/vendor/pdfjs/cmaps/';       //    pdfjsLib.workerSrc = 'js/vendor/pdf.worker.js';        //this.pdfToText = function(buf) {       //console.log(file.path);       //console.log(ab2str(buf));       //console.log(new Buffer(ab2str(buf), 'binary'));       //const enc = new FileReader();       //const enc = new TextDecoder();       //console.log(ab2str(buf));      //}     //  return buf;     //  }     //    bufView[i] = str.charCodeAt(i);     //  for (var i=0, strLen=str.length; i < strLen; i++) {     //  var bufView = new Uint16Array(buf);       //var buf = new ArrayBuffer(str.length*2); // 2 bytes for each char     //function str2ab(str) {        //console.log(buf.toString('utf-8'));       //}       //});       //  console.log(data);       //  if (err) return console.log(err);       //pdfExtract.extract(arr, options, (err,data) => {       //const options = {};       //const pdfExtract = new PDFExtract();       //})       //  console.log(data.text);       //pdf().then(function(data) {       //}); ad  F   �     ]   �  �  �  r  e  X  N  ,  
  �  �  �  w  9  �  �  �  �  �  �  �  �  �  �  �  �  }  Y  1    �  �  �  s  �
  =
  �	  	  �  �  u  B    �  �  �  �  _  ;  ~  _  ^  Z  V  U  9  4  0  /    �  �  �  �  �  �  {  p  h  d  c  b  H  4      �  �  ,    �  �  �  ]     �  B  �  �  �  �  �  �  �                                                                        }            }         };           }             myAudioItems.childNodes[this.state.indexAudioElement].play();             const indexAudioElement = Array.prototype.indexOf.call(myAudioItems.children, event.currentTarget) + 1;             const myAudioItems = document.getElementById('myAudioFiles');           if (allAudioElements && allAudioElements.length && allAudioElements.length >= 2) {           //allAudioElements[0].remove();            console.log(event.currentTarget);           const allAudioElements = audioTagName;         el.onended = (event) => {       for (let el of audioTagName) {     if (document.getElementById('playAllTheWords').checked && audioTagName && audioTagName.length && !Object.keys(audioTagName)[0].onended) {     const audioTagName = document.getElementsByTagName('audio');     });         event.target.value       noDatabaseFile:     this.setState({   checkBox = (event) => {     }     });         ''       textareaIsEmpty:     this.setState({     });         event.target.value       value:     this.setState({     console.log(this.state.value);   handleTextChange = (event) => {    }        previewFile = (file) => {    } 		}  			reader.readAsDataURL(file); 			reader.onload = (function(aImg) { return function(e) { aImg.src = e.target.wordIdItems; }; })(img); //if the file is an image, insert the content of the imageas the image in the dropbox 			const reader = new FileReader(); 			preview.appendChild(document.createElement('br'));                          //===END FILE PREVIEW AFTER DROP==// 			preview.appendChild(fileName); 			fileName.target = "_blank"; 			fileName.href = URL.createObjectURL(file); 			fileName.textContent = file.name+ ' (preview)';                         fileName.className += '.obj'; 			const fileName = document.createElement('a');                         //===FILE PREVIEW AFTER DROP==// 			if(file.type===('')) { preview.appendChild(noFileType); } // Assuming that "preview" is the div output where the content will be displayed. 			if(file.type.startsWith('text/')) { preview.appendChild(myImage); } // Assuming that "preview" is the div output where the content will be displayed. 			if(file.type.startsWith('application/')) { preview.appendChild(myImage); } // Assuming that "preview" is the div output where the content will be displayed. 			if(file.type.startsWith('image/')) { preview.appendChild(img); } // Assuming that "preview" is the div output where the content will be displayed. 			const preview = document.getElementById("preview");                         img.width = 60;                         img.height = 60; 			img.file = file; 			noFileType.src = `notype.png`; 			const noFileType = new Image(60,60); 			myImage.src = `application.png`; 			const myImage = new Image(60,60); 			img.classList.add("obj"); 			const img = document.createElement("img"); 			if (!file.type.startsWith('image/') && !file.type.startsWith('application/') && !file.type.startsWith('text/') && !file.type ===('')){ continue } 			const file = files[i]; 		for (let i = 0; i < files.length; i++) {   dropbox = (files) => {    }      //});     //  }     //    (rows[item.y] = rows[item.y] || []).push(item.text);     //    // accumulate text items into rows object, per line     //  } else if (item.text) {     //    rows = {}; // clear rows for next page     //    console.log("PAGE:", item.page);     //    printRows();     //    // end of file, or page     //  if (!item || item.page) {     //) {     //  item     //  err,     //new pdfreader.PdfReader().parseFileItems(file, function(     //     //}     //    .forEach(y => console.log((rows[y] || []).join(""))); 